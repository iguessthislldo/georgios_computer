module alu(r, op, A, B)
    input op
endmodule
