module alu(r, op, a, b)
    output [0:7] r;
    input op;
    input [0:7] a, b;
endmodule
