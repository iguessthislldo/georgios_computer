module mux(out, select, a, b);
    input select, a, b;
    output out;
endmodule
